* C:\Users\DELL\eSim-Workspace\MOD-10_Ripple\MOD-10_Ripple.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/08/22 20:29:45

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
scmode1  SKY130mode		
U3  clkIN rst Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
v4  rst GND pulse		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ mod_10		
U5  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ q1 q2 q3 q4 dac_bridge_4		
U4  q1 plot_v1		
U7  q2 plot_v1		
U8  q3 plot_v1		
U6  q4 plot_v1		
U9  rst plot_v1		
X1  vd vs Net-_SC3-Pad2_ Net-_SC1-Pad1_ clkIN GND avsd_opamp		
SC2  Net-_SC1-Pad1_ clkIN VDD sky130_fd_pr__res_generic_pd		
SC3  clkIN Net-_SC3-Pad2_ VDD sky130_fd_pr__res_generic_pd		
SC4  Net-_SC3-Pad2_ GND VDD sky130_fd_pr__res_generic_pd		
SC1  Net-_SC1-Pad1_ GND sky130_fd_pr__cap_mim_m3_1		
v1  vd GND DC		
U1  clkIN plot_v1		
v2  VDD GND DC		
v3  vs GND DC		

.end
